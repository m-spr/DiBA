------ ****  MAP4 with RECURSION  ***** --------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.All;

ENTITY MAPn_recursion IS 
  GENERIC(
	  h : INTEGER := 3;
	  a : INTEGER := 5;
	  b : INTEGER := 4;
	  c : INTEGER := 3;
	  d : INTEGER := 1;
	  e : INTEGER := 1;
	  f : INTEGER := 1;
	  k : INTEGER := 4 ---n0
		);
  PORT (clk,  rst,  run,  pause : IN STD_LOGIC ;
      reg_out : OUT STD_LOGIC;
	  din : IN STD_LOGIC_VECTOR(16*a*b*c*d*e*f -1 DOWNTO 0);
	  w : IN STD_LOGIC_VECTOR(16*a*b*c*d*e*f -1 DOWNTO 0);
	  dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
		  );
END MAPn_recursion;	  



ARCHITECTURE behavioral_MAPn OF MAPn_recursion IS 


COMPONENT MAPn_recursion IS 
  GENERIC(
	  h : INTEGER := 3;
	  a : INTEGER := 5;
	  b : INTEGER := 4;
	  c : INTEGER := 3;
	  d : INTEGER := 1;
	  e : INTEGER := 1;
	  f : INTEGER := 1;
	  k : INTEGER := 4 ---n0
		);
  PORT (clk,  rst,  run,  pause : IN STD_LOGIC ;
      reg_out : OUT STD_LOGIC;
	  din : IN STD_LOGIC_VECTOR(16*a*b*c*d*e*f -1 DOWNTO 0);
	  w : IN STD_LOGIC_VECTOR(16*a*b*c*d*e*f -1 DOWNTO 0);
	  dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
		  );
END COMPONENT;
		
COMPONENT  MAP_1 IS 
GENERIC(
      n : INTEGER := 15
        );
PORT ( 
      clk,  rst ,add_reg , reg_out: IN STD_LOGIC;
      din : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
      w : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
      dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	   );

END COMPONENT;

COMPONENT CAP IS 
  GENERIC(
      n : INTEGER := 16
        );
  PORT ( clk, rst, run : IN STD_LOGIC ;
        reg_OUT : OUT STD_LOGIC;
	dIN : IN STD_LOGIC_VECTOR(32*n-1 DOWNTO 0);
        dout: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
       );
END COMPONENT;

SIGNAL rego : STD_LOGIC_VECTOR (a DOWNTO 1 );
SIGNAL regocap , wait_data_out: STD_LOGIC_VECTOR (h+1 DOWNTO 0 ) := (others => '0');
	

SIGNAL data_out_map : STD_LOGIC_VECTOR(32*a -1 DOWNTO 0);
	
BEGIN 

	regocap(h) <= run;

			h0 : if h = 1 generate
				MAP_1s: FOR I IN 1 TO a GENERATE
		    MAP1 :  MAP_1
		        GENERIC MAP( k )
				PORT MAP (  
			        clk,  rst,  run,  rego(I),
				din(((I*16)-1) DOWNTO ((I-1)*16)),  
				w(((I*16)-1) DOWNTO ((I-1)*16)),  
				data_out_map((I*32)-1 DOWNTO (I-1)*32)
						);
				END GENERATE MAP_1s;
			CAP_1 : CAP 
				GENERIC MAP (a)
					PORT MAP( 
						clk,  rst,  rego(1),  
						regocap(0),  
						data_out_map,  
						dout
						);
			end generate h0;
			
			hb0 : if h > 1 generate
				MAP_ns_for : FOR i in 1 to a generate
			MAP_ns : MAPn_recursion 
			    GENERIC map( h-1, b, c, d, e, f, 1, k )
				    PORT map(clk,  rst,  regocap(h),  pause,
						rego(i), 
						din (16*b*c*d*e*f*(i) -1 downto 16*b*c*d*e*f*(i-1)),
						w (16*b*c*d*e*f*(i) -1 downto 16*b*c*d*e*f*(i-1)),
						data_out_map((32*i)-1 downto 32*(i-1)) 
					     );   
				END GENERATE MAP_ns_for;
			CAP_n : CAP 
				GENERIC MAP (a)
					PORT MAP( 
						clk,  rst,  rego(1),  
						regocap(h-1),
						data_out_map,  
						dout
					     );
			END GENERATE hb0;
				
				
	reg_out <= regocap(h-1);
END behavioral_MAPn;



--------------------------------------------------------------
LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY MAPn_tb IS

END MAPn_tb;	  

ARCHITECTURE tb OF MAPn_tb Is

Component MAPn_recursion IS 
  GENERIC(
	  h : INTEGER := 2;
	  a : INTEGER := 5;
	  b : INTEGER := 4;
	  c : INTEGER := 3;
	  d : INTEGER := 1;
	  e : INTEGER := 1;
	  f : INTEGER := 1;
	  k : INTEGER := 4 ---n0
		);
  PORT (clk,  rst,  run,  paUSE : IN STD_LOGIC ;
      reg_OUT : OUT STD_LOGIC;
	  din : IN STD_LOGIC_VECTOR(16*a*b*c*d*e*f -1 DOWNTO 0);
	  w : IN STD_LOGIC_VECTOR(16*a*b*c*d*e*f -1 DOWNTO 0);
	  dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
		  );  
END COMPONENT;

SIGNAL clk, rst, run, paUSE :  STD_LOGIC := '1';
SIGNAL reg_OUT : STD_LOGIC ;
SIGNAL din : STD_LOGIC_VECTOR(16*5*4*3*1*1*1 -1 DOWNTO 0);
SIGNAL w : STD_LOGIC_VECTOR(16*5*4*3*1*1*1 -1 DOWNTO 0);
SIGNAL dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
		
BEGIN 

MAPn : MAPn_recursion  
  GENERIC MAP(3, 3, 4, 5, 1, 1, 1, 7)
  PORT MAP (clk,  rst,  run,  paUSE,
      reg_OUT ,
	  din , w ,
	  dout  ); 
		  
clk <= not clk AFTER 5 ns;
rst <= '0' AFTER 30 ns;
run <= '0',  '1' AFTER 50 ns;
paUSE <= '0'; -- , '1' AFTER 180 ns , '0' AFTER 200 ns, '1' AFTER 480 ns , '0' AFTER 600 ns;
din <= "000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001";
w <= "000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001";
END tb;



